library verilog;
use verilog.vl_types.all;
entity somador4_vlg_vec_tst is
end somador4_vlg_vec_tst;
