library verilog;
use verilog.vl_types.all;
entity cod_hamming_vlg_vec_tst is
end cod_hamming_vlg_vec_tst;
