library verilog;
use verilog.vl_types.all;
entity injeta_erro_vlg_vec_tst is
end injeta_erro_vlg_vec_tst;
