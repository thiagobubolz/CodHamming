library verilog;
use verilog.vl_types.all;
entity decod_hamming_vlg_vec_tst is
end decod_hamming_vlg_vec_tst;
